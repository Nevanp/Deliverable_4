module channel(
    input clk,
    input signed [17:0] x_in,
    output reg signed [17:0] y
);


endmodule