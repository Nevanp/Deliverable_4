module upconv(
    input clk,
    input sym_clk,
    input sam_clk,
    input signed [17:0] x_in,
    output reg signed [17:0] y
);

endmodule